`include "cpu_defs.svh"

module trivial_mips(
	input  clk, rst,
	input  WishboneReq_t ibus_i,
	output WishboneRes_t ibus_o,
	input  WishboneReq_t dbus_i,
	output WishboneRes_t dbus_o
);


endmodule

module ctrl(
	input rst,
	input stall_from_id,
	input stall_from_ex,
	input stall_from_mem,
	input stall_from_wb
);

endmodule

`ifndef COMMON_DEFS_SVH
`define COMMON_DEFS_SVH

/*
    Options to control functional parts to be compiled
*/

`define ENABLE_CPU_FPU                  1
`define ENABLE_PERIPHERAL_ETHERNET      1
`define ENABLE_PERIPHERAL_FLASH         1
`define ENABLE_PERIPHERAL_GPIO          1
`define ENABLE_PERIPHERAL_GRAPHICS      1
`define ENABLE_PERIPHERAL_TIMER         1
`define ENABLE_PERIPHERAL_UART          1
`define ENABLE_PERIPHERAL_USB           1

`endif
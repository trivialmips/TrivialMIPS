`include "common_defs.svh"

module sram_controller(
    Bus_if.slave   inst_bus,
    Bus_if.salve   data_bus,
    Sram_if.master base_ram,
    Sram_if.master ext_ram
);


endmodule
`include "cpu_defs.svh"

module reg_pc(
	input  clk, rst,
	output ce,   // chip enable
	output InstAddr_t addr
);

endmodule
